
`include "timescale.v"

// synthesis attribute priority_extract of count_leading_zeroes is force

module count_leading_zeroes(
	in,

	count
);

input	[30:0]	in;

output	[4:0]	count;

reg	[4:0]	count;


always @(in)
begin
	// The if/else form is recommended by the Xilinx XST user's guide
	// for inferring a priority encoder:
	if      (in[30])	count = 5'h0;
	else if (in[29])	count = 5'h1;
	else if (in[28])	count = 5'h2;
	else if (in[27])	count = 5'h3;
	else if (in[26])	count = 5'h4;
	else if (in[25])	count = 5'h5;
	else if (in[24])	count = 5'h6;
	else if (in[23])	count = 5'h7;
	else if (in[22])	count = 5'h8;
	else if (in[21])	count = 5'h9;
	else if (in[20])	count = 5'ha;
	else if (in[19])	count = 5'hb;
	else if (in[18])	count = 5'hc;
	else if (in[17])	count = 5'hd;
	else if (in[16])	count = 5'he;
	else if (in[15])	count = 5'hf;
	else if (in[14])	count = 5'h10;
	else if (in[13])	count = 5'h11;
	else if (in[12])	count = 5'h12;
	else if (in[11])	count = 5'h13;
	else if (in[10])	count = 5'h14;
	else if (in[9])		count = 5'h15;
	else if (in[8])		count = 5'h16;
	else if (in[7])		count = 5'h17;
	else if (in[6])		count = 5'h18;
	else if (in[5])		count = 5'h19;
	else if (in[4])		count = 5'h1a;
	else if (in[3])		count = 5'h1b;
	else if (in[2])		count = 5'h1c;
	else if (in[1])		count = 5'h1d;
	else if (in[0])		count = 5'h1e;
	else			count = 5'hx;

/*
	casez(in)
	31'b1??????????????????????????????: count = 5'h0;
	31'b01?????????????????????????????: count = 5'h1;
	31'b001????????????????????????????: count = 5'h2;
	31'b0001???????????????????????????: count = 5'h3;
	31'b00001??????????????????????????: count = 5'h4;
	31'b000001?????????????????????????: count = 5'h5;
	31'b0000001????????????????????????: count = 5'h6;
	31'b00000001???????????????????????: count = 5'h7;
	31'b000000001??????????????????????: count = 5'h8;
	31'b0000000001?????????????????????: count = 5'h9;
	31'b00000000001????????????????????: count = 5'ha;
	31'b000000000001???????????????????: count = 5'hb;
	31'b0000000000001??????????????????: count = 5'hc;
	31'b00000000000001?????????????????: count = 5'hd;
	31'b000000000000001????????????????: count = 5'he;
	31'b0000000000000001???????????????: count = 5'hf;
	31'b00000000000000001??????????????: count = 5'h10;
	31'b000000000000000001?????????????: count = 5'h11;
	31'b0000000000000000001????????????: count = 5'h12;
	31'b00000000000000000001???????????: count = 5'h13;
	31'b000000000000000000001??????????: count = 5'h14;
	31'b0000000000000000000001?????????: count = 5'h15;
	31'b00000000000000000000001????????: count = 5'h16;
	31'b000000000000000000000001???????: count = 5'h17;
	31'b0000000000000000000000001??????: count = 5'h18;
	31'b00000000000000000000000001?????: count = 5'h19;
	31'b000000000000000000000000001????: count = 5'h1a;
	31'b0000000000000000000000000001???: count = 5'h1b;
	31'b00000000000000000000000000001??: count = 5'h1c;
	31'b000000000000000000000000000001?: count = 5'h1d;
	31'b0000000000000000000000000000001: count = 5'h1e;
	default: count = 5'h0;
	endcase
*/
end

endmodule
